library ieee;
use ieee.std_logic_1164.all;

entity rom_cm is
    generic(n : integer := 64);
    port(
        a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12 : out std_logic_vector(n-1 downto 0)
    );
end;

architecture arch of rom_cm is
begin
    a1 <= "1111011001100110011001100110011001100110011001100110011010000000"; ---0.60
    a2 <= "1111111001100110011001100110011001100110011001100110011001100000"; ---0.10
    a3 <= "0001000110011001100110011001100110011001100110011001101000000000"; -- 1.10
    a4 <= "0000001100110011001100110011001100110011001100110011001101000000"; -- 0.20
    a5 <= "1111001100110011001100110011001100110011001100110011001100000000"; ---0.80
    a6 <= "0000100110011001100110011001100110011001100110011001100110000000"; -- 0.60
    a7 <= "1111010011001100110011001100110011001100110011001100110100000000"; ---0.70
    a8 <= "0000101100110011001100110011001100110011001100110011001100000000"; -- 0.70
    a9 <= "0000101100110011001100110011001100110011001100110011001100000000"; -- 0.70
    a10 <= "0000010011001100110011001100110011001100110011001100110011000000"; -- 0.30
    a11 <= "0000100110011001100110011001100110011001100110011001100110000000"; -- 0.60
    a12 <= "0000111001100110011001100110011001100110011001100110011010000000"; -- 0.90
end;
