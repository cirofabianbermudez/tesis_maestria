LIBRARY UNISIM;
USE UNISIM.vcomponents.ALL;
